// Module - Sync Unit Ouput Module 
// Author: James Ashie Kotey
// Adapted from hv_sync_generator by Urish - VGA-Playground.com 

/*
    Description: 
        Generates sync pulses for VGA monitor, (H-SYNC ,V-SYNC) targeted to 640 * 480 output, 
        Pixel coordinates for the graphics controller,§
        and sync signals for the game logic units.  
*/

module sync_generator (  
    input              clk,
    input              reset,
    output reg         hsync,
    output reg         vsync,
    output wire        display_on,
    output wire [9:0]  screen_hpos,
    output wire [9:0]  screen_vpos,
    output wire        frame_end,
    output wire        input_enable
);
    
    reg [9:0] hpos = 0;
    reg [9:0] vpos = 0;

    // declarations for TV-simulator sync parameters

    // horizontal constants

    parameter H_DISPLAY = 640;  // horizontal display width
    parameter H_BACK = 48;  // horizontal left border (back porch)
    parameter H_FRONT = 16;  // horizontal right border (front porch)
    parameter H_SYNC = 96;  // horizontal sync width

    // vertical constants

    parameter V_DISPLAY = 480;  // vertical display height
    parameter V_TOP = 33;  // vertical top border
    parameter V_BOTTOM = 10;  // vertical bottom border
    parameter V_SYNC = 2;  // vertical sync # lines

    // derived constants

    parameter H_SYNC_START = H_DISPLAY + H_FRONT;
    parameter H_SYNC_END = H_DISPLAY + H_FRONT + H_SYNC - 1;
    parameter H_MAX = H_DISPLAY + H_BACK + H_FRONT + H_SYNC - 1;
    parameter V_SYNC_START = V_DISPLAY + V_BOTTOM;
    parameter V_SYNC_END = V_DISPLAY + V_BOTTOM + V_SYNC - 1;
    parameter V_MAX = V_DISPLAY + V_TOP + V_BOTTOM + V_SYNC - 1;

    wire hmaxxed = (hpos == H_MAX) || reset;  // set when hpos is maximum
    wire vmaxxed = (vpos == V_MAX) || reset;  // set when vpos is maximum
    
    wire hblanked = (hpos == H_DISPLAY);
    wire vblanked = (vpos == V_DISPLAY);

    assign screen_hpos = (hpos < H_DISPLAY)? hpos : 0; 
    assign screen_vpos = (vpos < V_DISPLAY)? vpos : 0;

    // horizontal position counter

    always @(posedge clk) begin

        if (reset) begin
            hpos <= 0;
            hsync <= 0; // active high pulse
        end 

        else begin
            hsync <= (hpos >= H_SYNC_START && hpos <= H_SYNC_END);
            if (hmaxxed) begin
            hpos <= 0;
            end else begin
            hpos <= hpos + 1;
            end
        end
    end

    // vertical position counter

    always @(posedge clk) begin

        if (reset) begin
            vpos <= 0;
            vsync <= 0;  // active high pulse
        end
        
        else begin
            vsync <= (vpos >= V_SYNC_START && vpos <= V_SYNC_END);
            if (hmaxxed)
            if (vmaxxed) begin
            vpos <= 0;
            end else begin
                vpos <= vpos + 1;
            end
        end
    end

    // display_on is set when beam is in "safe" visible frame
    assign display_on = (hpos < H_DISPLAY) && (vpos < V_DISPLAY);
    assign frame_end = hblanked && vblanked;
    assign input_enable = 1; //(hblanked && vpos < V_DISPLAY);

endmodule
